/** Copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_clocking.cdl
 * @brief Testbench for numerous clocking modules
 *
 */
/*a Includes */
include "std::bit_delay.h"
include "clocking.h"
include "clocking_modules.h"

/*a Module */
module tb_clocking( clock clk,
                    input bit reset_n,
                    output t_bit_delay_config   delay_config_cpm,
                    output t_bit_delay_config   delay_config_cet,
                    input  t_bit_delay_response delay_response,
                    input  t_phase_measure_request measure_request,
                    output t_phase_measure_response measure_response,
                    input  t_eye_track_request eye_track_request,
                    output t_eye_track_response  eye_track_response,
                    input  bit[4] data_p_in,
                    input  bit[4] data_n_in
)
{

    /*b Nets */
    net t_bit_delay_config   delay_config_cpm;
    net t_bit_delay_config   delay_config_cet;
    // net t_bit_delay_response delay_response;
    // net t_phase_measure_request measure_request;
    net t_phase_measure_response measure_response;
    // net t_eye_track_request  eye_track_request;
    net t_eye_track_response eye_track_response;
    // net bit[4] data_p_in;
    // net bit[4] data_n_in;

    /*b Instantiations */
    instantiations: {
        clocking_phase_measure cpm(clk <- clk,
                                   reset_n <= reset_n,
                                   delay_config   => delay_config_cpm,
                                   delay_response <= delay_response,
                                   measure_request <= measure_request,
                                   measure_response => measure_response );
        clocking_eye_tracking cet(clk <- clk,
                                  data_clk <- clk,
                                  reset_n <= reset_n,
                                  data_p_in <= data_p_in,
                                  data_n_in <= data_n_in,
                                  delay_config   => delay_config_cet,
                                  delay_response <= delay_response,
                                  eye_track_request <= eye_track_request,
                                  eye_track_response => eye_track_response );
    }

    /*b All done */
}
