/** @copyright (C) 2016-2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   timer.cdl
 * @brief  Standardized 64-bit timer with synchronous control
 *
 * CDL implementation of a standard 64-bit timer using synchronous control.
 *
 */
/*a Constants */
/*v sync_toggle_count
 *
 * This is the number of toggle cycles to operate on for counting
 *  early/late/unexpected toggles.
 * A toggle cycle is indicated by the master time value crossing the
 * first-to-second quarter-window boundary.
 * If this occurs when the slave timer value is still in the first
 * quarter window then the slave is deemed late
 * If this occurs when the slave timer value is still in the second
 * quarter window then the slave is deemed early
 * If this occurs in the other half of the window we have an unexpected
 * value - and this causes the system to be marked as out of lock.
 *
 * The maximum retard/advance is once per this number of toggles
 *
 * The time between retard/advances is then once per:
 *    sync_toggle_count * toggle_period 
 *
 * The standard timer adjusts by 1/2 a slave clock tick per retard/advance
 *
 * For a 100MHz slave (10ns clock period) the retard/advance adjustment is 5ns.
 * For sync_toggle_count of 16 with toggle_period of 512ns (i.e ~8200 ns) this
 * accounts for 600ppm
 *
 * For a 600MHz slave (1.6ns clock period) the retard/advance adjustment is 800ps.
 * For sync_toggle_count of 16 with toggle_period of 256ns (i.e ~4000 ns) this
 * accounts for 200ppm
 *
 * Note that the ppm here should be the sum of all clocks and long-term PLL jitter
 * leading to the slave clock
 *
 * T.period(ns)  STC  AdjPeriod Clk(MHz) Clk(ns)  Adj(ns)  ppm
 *    64         16     1.0us     1000     1.0       0.5   488
 *    64         16     1.0us      600     1.6       0.8   780
 *    64         16     1.0us      500     2.0       1.0   977
 *    64         16     1.0us      250     4.0       2.0  1954
 *
 *   128         16     2.0us     1000     1.0       0.5   244
 *   128         16     2.0us      600     1.6       0.8   390
 *   128         16     2.0us      500     2.0       1.0   488
 *   128         16     2.0us      250     4.0       2.0   977
 *   128         16     2.0us      125     8.0       4.0  1954
 *
 *   256         16     4.1us     1000     1.0       0.5   122
 *   256         16     4.1us      600     1.6       0.8   195
 *   256         16     4.1us      500     2.0       1.0   244
 *   256         16     4.1us      250     4.0       2.0   488
 *   256         16     4.1us      125     8.0       4.0   976
 *   256         16     4.1us       64    15.6       7.8  1906
 *
 *   512         16     8.2us     1000     1.0       0.5    61
 *   512         16     8.2us      600     1.6       0.8    98
 *   512         16     8.2us      500     2.0       1.0   122
 *   512         16     8.2us      250     4.0       2.0   244
 *   512         16     8.2us      125     8.0       4.0   488
 *   512         16     8.2us       64    15.6       7.8   953
 *
 *  1024         16    16.4us      500     2.0       1.0    61
 *  1024         16    16.4us      250     4.0       2.0   122
 *  1024         16    16.4us      125     8.0       4.0   244
 *  1024         16    16.4us       64    15.6       7.8   477
 *  1024         16    16.4us       32    31.2      15.6   954
 *
 *  2048         16    32.8us      250     4.0       2.0    61
 *  2048         16    32.8us      125     8.0       4.0   122
 *  2048         16    32.8us       64    15.6       7.8   238
 *  2048         16    32.8us       32    31.2      15.6   477
 *
 *  4096         16    65.5us      125     8.0       4.0    61
 *  4096         16    65.5us       64    15.6       7.8   119
 *  4096         16    65.5us       32    31.2      15.6   238
 *  4096         16    65.5us       10   100.0      50.0   763
 *
 * Table shows ppm of >50 and T.period>=16 clock periods
 *
 * AdjPeriod is T.period * STC
 *
 * Clock period is 1000.0 / Clk(MHz)
 *
 * The adjustment is half the clock period
 *
 * The ppm is adjustment / AdjPeriod
 *
 * To support the range of clocks from 10MHz to 1GHz a selection of
 *  64ns, 256ns, 1024ns and 4096ns seems sensible
 * This corresponds to LSB of 4, 6, 8 and 10 for the quater-window size
 *
 * LSB of 4 (period 64ns) should be used for clocks of >=250MHz
 * LSB of 6 (period 256ns) should be used for clocks of 64MHz to 250MHz
 * LSB of 8 (period 1us) should be used for clocks of 32MHz to 64MHz
 * LSB of 10 (period 4us) should be used for clocks of 8MHz to 32MHz
 *
 */
constant integer sync_toggle_count=16;
constant integer toggle_count_width = sizeof(2*sync_toggle_count-1);

/*a Includes
 */
include "std::tech_sync.h"
include "clock_timer.h"
include "clock_timer_modules.h"

/*a Types */
/*t t_slave_fsm
 *
 * State of the slave timer FSM, in the slave clock domain
 *
 */
typedef fsm {
    slave_fsm_idle                {
        slave_fsm_toggle_complete
    } "Waiting for master toggle to be detected";
    slave_fsm_toggle_complete     {
        slave_fsm_idle
    } "Recorded toggle, if last toggle of window then update timer; go back to idle";
} t_slave_fsm;

/*t t_slave_action
 *
 * Transition that the slave FSM and state needs to perform in this slave clock cycle
 *
 */
typedef enum [4] {
    slave_action_none                "No toggle seen, nothing to do",
    slave_action_idle                "Return to idle (from @a toggle_complete)",
    slave_action_simultaneous_toggle "Master toggle detected at same time as slave timer value crossed window",
    slave_action_slave_early         "Master toggle detected while slave timer value is already in second quarter",
    slave_action_slave_late          "Master toggle detected while slave timer value is still in first quarter",
    slave_action_unexpected_toggle   "Master toggle detected while slave timer value is way off",
    slave_action_not_locked          "Mark as not locked and return to idle",
    slave_action_locked              "Mark as locked with no need to change slave timer value and return to idle",
    slave_action_locked_retard       "Mark as locked with slave timer ahead (hence request slave timer retard) and return to idle",
    slave_action_locked_advance      "Mark as locked with slave timer behing (hence request slave timer advance) and return to idle",
} t_slave_action;

/*t t_timing_op
 *
 * Enumeration of timer operations that can be performed - nothing, advance or retard
 *
 */
typedef enum [2] {
    timing_op_none,
    timing_op_advance,
    timing_op_retard
} t_timing_op;

/*t t_slave_combs
 *
 * Combinatorial decode of the slave state
 *
 */
typedef struct {
    bit     master_toggle      "Asserted if the slave has seen the master cross the quarter-window boundary";
    bit[64] top_value          "Top bits of timer value, bottom window_bits downward zeroed out";
    bit     top_value_matches  "Asserted if master and slave timer values through the mask are equal - if this is not the case on a toggle then there is no lock";
    bit[2]  window_bits        "Selected slave timer value bits for the quarter window";
    t_slave_action action      "Action for the slave state machine";
    bit[toggle_count_width] toggle_diff "Difference in early and late toggle counts for the slave in the current set of toggles";
    bit toggles_close_enough            "Valid after enough toggles seen, asserted if the slave timer value has crosssed the window nearly as often early as late (and vice versa)";
    bit more_early_toggles              "Asserted if the slave timer value has crossed the window early more than late";
} t_slave_combs;

/*t t_slave_toggles
 *
 * State in the slave that counts the toggles
 *
 */
typedef struct {
    bit[toggle_count_width] seen        "Count of master quarter-window crossing seen";
    bit[toggle_count_width] early       "Number of times the slave was early within @a seen";
    bit[toggle_count_width] late        "Number of times the slave was late within @a seen";
    bit                     unexpected  "Set if the slave was ever late within @a seen";
} t_slave_toggles;

/*t t_slave_window
 *
 * State about the slave timer value, used to determine if the slave timer value is on time, late or early
 *
 */
typedef struct {
    bit value_in_first_quarter   "Asserted if in the first quarter of the timer value window (window bits are 2b00)";
    bit value_in_second_quarter  "Asserted if in the second quarter of the timer value window (window bits are 2b01)";
} t_slave_window;

/*t t_slave_state
 *
 */
typedef struct {
    bit last_master_quarter_window_passed   "Used for edge detection on sync version of quarter_window_passed";
    bit[2] last_window_bits                 "The quarter-window bits of the slave time value in the last slave clock tick";
    t_slave_window window                   "Which quarter-window the slave timer value is in - first, second, or neither";
    t_slave_window last_window              "Which quarter-window the slave timer value was in during the last cycle";
    t_slave_window ancient_window           "Which quarter-window the slave timer value was in during the last cycle but one";
    t_slave_fsm fsm_state                   "Slave FSM state";
    t_slave_toggles toggles                 "Toggle counts for the slave FSM";
    bit synchronize_request                 "Slave clock record of the synchronized master 'synchronize' request going high - used to determine if synchronization is required";
    t_timing_op request_timing              "Request to timer control to advance/retard - but only if locking enabled";
    t_timer_control timer_control           "Timer control to the internal slave clock_timer and for the @a slave_timer_control_out";
    bit phase_locked                        "Asserted if phase locked to master";
    bit locked                              "Asserted if phase locked to master and upper value bits match";
} t_slave_state;

/*t t_master_combs
 *
 * Combinatorial decode of the master side - some also used for the slave side if the input controls are 'configuration' slow
 *
 */
typedef struct {
    bit[64] top_value_mask  "Mask of top bits of timer value dependent on input control window size - used by master and slave";
    bit[64] quarter_window  "Bits 01 in the quarter-window position - just below top_value_mask - used by master and slave";
    bit[64] top_value       "Top bits of timer value, bottom window_bits downward zeroed out - used by master, and by slave just after end of first quarter window";
    bit[2]  window_bits     "Two bits of timer value indicate which quarter window it is in";
} t_master_combs;

/*t t_master_state
 *
 */
typedef struct {
    bit synchronize_pending    "Asserted if master timer control has synchronize set at some point, until request is taken";
    bit synchronize_request    "Asserted if @a synchronize_pending was asserted when the first quarter window was passed (so @a top_value will be stable for slave clock); high for a whole window";
    bit quarter_window_passed  "Asserted when the quarter window is passed";
    bit[2] last_window_bits    "Last value of first 2 bits of window";
} t_master_state;

/*a Module */
module clock_timer_async( clock master_clk             "Master clock",
                          input bit master_reset_n     "Active low reset",
                          clock slave_clk              "Slave clock, asynchronous to master",
                          input bit slave_reset_n     " Active low reset",
                          input t_timer_control  master_timer_control     "Timer control in the master domain - synchronize, reset, enable and lock_to_master are used",
                          input t_timer_value    master_timer_value       "Timer value in the master domain - only 'value' is used",
                          input t_timer_control   slave_timer_control_in  "Timer control in the slave domain - only adder values are used",
                          output t_timer_control  slave_timer_control_out "Timer control in the slave domain for other synchronous clock_timers - all valid",
                          output t_timer_value    slave_timer_value       "Timer value in the slave domain"
    )
"""
Module to take a timer control in one clock domain and synchronize it to another clock domain.

It operates using a window in the timer values, that starts at a particular (run time) bit of the timer value.
This window is separated into four quarters.
For example, the window boundary can be at intervals of 1024; hence quarter windows are at intervals of 256.
The timer value is in the first quarter if, modulo 1024, its value is 0 to 255. It is in the second quarter 
if, modulo 1024, its value is 256 to 511.

The module uses the crossing from the first quarter to the second quarter as a 'toggle'. At this point,
given suitable configuration of the window size, the slave is guaranteed to see the top (non window) bits of
the master time value as stable.

The slave should also see its timer value cross the quarter window in the same slave clock tick as it sees the master
timer value cross the quarter window. The phase difference between when these toggles occur can be used to
advance or retard the slave clock.

The slave has to operate on synchronized versions of the master toggle, and this takes a couple of slave
clock ticks to stabilize; hence the slave has to delay its slave timer value quarter window crossing
to match.

The 'enable', 'reset' and 'lock_to_master' are simply synchronized across.
The 'synchronize' control requires a small state machine - when this is asserted the master_timer_value
is monitored and when it crosses from quarter window boundary a control is passed to the
slave to inform it to synchronize to the upper master_timer_value bits at half the window size.
It is the rising edge of the synchronized signal (that must clearly occur only when the master timer value upper
bits are stable) that is used by the slave to invoke a synchronization (and storage of the master time value upper bits).
The lower bits of the slave timer can be set to the quarter window boundary (it will be a couple of slave clock ticks
behind the master at this point, but further 'advance' of the clock should bring it in to phase).

The slave monitors a synchronized version of the master toggle (master timer value crossing the quarter window boundary).
If this occurs when the slave has also just crossed the boundary then the toggle is deemed 'simultaneous'.
If the master crosses while the slave is still in the first quarter, then the slave is late.
If the master crosses when the slave had already moved into the second quarter, then the slave was early.
If the master crosses when the slave was in the third or fourth quarters then the slave is just out of lock.

A running count of early, late toggles and unexpected toggles is maintained.
After a number of master window crossings are seen the slave can retard or advance its clock, or report out of lock.
The counts are reset.
If more than one unexpected toggled occurs then the timer is deemed 'not locked'.
"""
{
    /*b Master state */
    default clock master_clk;
    default reset active_low master_reset_n;
    clocked t_master_state master_state= {*=0} "State of the master";
    comb    t_master_combs master_combs        "Combinatorial decode of the master";
    
    /*b Handle the master side */
    master_logic """
    The master side monitors the quarter window boundary, and toggles its @a quarter_window_passed state whenever the
    timer value crosses from the first quarter to the second quarter.

    It also maintains the synchronization request - it records if a synchronize is performed on the control in, and
    will change its @a synchronize_request signal on the quarter window boundary so that the slave can synchronize it,
    and use negative edge detection to determine a synchronization is required.
    """: {
       
        if (master_timer_control.synchronize!=0) {
            master_state.synchronize_pending <= 1;
        }
        master_state.last_window_bits <= master_combs.window_bits;
        if ((master_combs.window_bits==2b01) &&
            (master_state.last_window_bits==2b00)) {
            master_state.quarter_window_passed <= !master_state.quarter_window_passed;
            master_state.synchronize_request   <= 0;
            if (master_state.synchronize_pending && !master_state.synchronize_request) {
                master_state.synchronize_request <= 1;
                master_state.synchronize_pending <= 0;
            }
        }
    }

    /*b Synchronizers to slave */
    net bit slave_sync_master_reset_counter;
    net bit slave_sync_master_enable_counter;
    net bit slave_sync_master_lock_to_master;
    net bit slave_sync_master_synchronize_request;
    net bit slave_sync_master_quarter_window_passed;
    slave_synchronizers """
    Synchronization from the master to the slave domain.

    @a reset_counter, @a enable_counter and @a lock_to_master are slow and level sensitive

    @a synchronize_request is negative edge detected

    @a quarter_window_passed toggles and every edge is detected
    """: {
        tech_sync_bit slave_reset_counter_flop(clk <- slave_clk, reset_n<=slave_reset_n,
                                               d <= master_timer_control.reset_counter,
                                               q => slave_sync_master_reset_counter ); // level sensitive
        tech_sync_bit slave_enable_counter_flop(clk <- slave_clk, reset_n<=slave_reset_n,
                                               d <= master_timer_control.enable_counter,
                                               q => slave_sync_master_enable_counter ); // level sensitive
        tech_sync_bit slave_lock_to_master_flop(clk <- slave_clk, reset_n<=slave_reset_n,
                                               d <= master_timer_control.lock_to_master,
                                               q => slave_sync_master_lock_to_master ); // level sensitive
        tech_sync_bit slave_synchronize_flop(clk <- slave_clk, reset_n<=slave_reset_n,
                                             d <= master_state.synchronize_request,
                                             q => slave_sync_master_synchronize_request ); // rising edge important
        tech_sync_bit slave_window_flop(clk <- slave_clk, reset_n<=slave_reset_n,
                                        d <= master_state.quarter_window_passed,
                                        q => slave_sync_master_quarter_window_passed ); // toggle important
    }
    
    /*b Slave state */
    default clock slave_clk;
    default reset active_low slave_reset_n;
    clocked t_slave_state slave_state= {*=0} "State of the slave";
    comb    t_slave_combs slave_combs        "Combinatorial decode of slave state and controls";
    net     t_timer_value slave_timer_value  "Timer value from the slave clock domain clock_timer module";

    /*b Handle the slave side */
    slave_logic """
    """: {
        /*b Determine if top part (non window) of timer_value match between slave and master.
         *  This is only used at the quarter window boundary, and hence should be stable
         */
        slave_combs.top_value_matches = 0;
        if (master_combs.top_value==slave_combs.top_value) {
            slave_combs.top_value_matches = 1;
        }

        /*b Record quarter window bits for the slave, and history of
         *  which quarter the slave timer is in
         */
        slave_state.last_window_bits <= slave_combs.window_bits;
        slave_state.last_window      <= slave_state.window;
        slave_state.ancient_window   <= slave_state.last_window;
        if (slave_state.last_window_bits != slave_combs.window_bits) {
            slave_state.window.value_in_first_quarter   <= (slave_combs.window_bits==2b00);
            slave_state.window.value_in_second_quarter  <= (slave_combs.window_bits==2b01);
        }

        /*b Determine if master has toggled (hence crossed quarter
         *  window boundary), and calculate toggle count deltas and
         *  results
         */
        slave_state.last_master_quarter_window_passed <= slave_sync_master_quarter_window_passed;
        slave_combs.master_toggle = (slave_state.last_master_quarter_window_passed != slave_sync_master_quarter_window_passed);
        slave_combs.toggle_diff          = slave_state.toggles.early - slave_state.toggles.late;
        slave_combs.more_early_toggles   = slave_state.toggles.early > slave_state.toggles.late;
        slave_combs.toggles_close_enough = ( (slave_combs.toggle_diff[3;toggle_count_width-3]==0) ||
                                             (slave_combs.toggle_diff[3;toggle_count_width-3]==-1) );

        /*b Decode the slave FSM state and determine its action */
        slave_combs.action = slave_action_none;
        full_switch (slave_state.fsm_state) {
        case slave_fsm_idle: {
            if (slave_combs.master_toggle) {
                slave_combs.action = slave_action_unexpected_toggle;
                if (slave_state.last_window.value_in_first_quarter) {
                    slave_combs.action = slave_action_slave_late;
                } elsif (slave_state.last_window.value_in_second_quarter) {
                    if (slave_state.ancient_window.value_in_first_quarter) {
                        slave_combs.action = slave_action_simultaneous_toggle;
                    } else {
                      slave_combs.action = slave_action_slave_early;
                    }
                }
            }
        }
        case slave_fsm_toggle_complete: {
            if (slave_state.toggles.unexpected) {
                slave_combs.action = slave_action_not_locked;
            } elsif (slave_combs.toggles_close_enough) {
                slave_combs.action = slave_action_locked;
            } else {
                slave_combs.action = slave_action_locked_advance;
                if (slave_combs.more_early_toggles) {
                    slave_combs.action = slave_action_locked_retard;
                }
            }
            if (slave_state.toggles.seen != sync_toggle_count) {
                slave_combs.action = slave_action_idle;
            }
        }
        }

        /*b Perform the action required from the slave FSM state machine decode */
        full_switch (slave_combs.action) {
        case slave_action_none: {
            slave_state.fsm_state <= slave_state.fsm_state;
        }
        case slave_action_idle: {
            slave_state.fsm_state <= slave_fsm_idle;
        }
        case slave_action_simultaneous_toggle: {
            slave_state.fsm_state    <= slave_fsm_toggle_complete;
            slave_state.toggles.seen  <= slave_state.toggles.seen + 1;
        }
        case slave_action_slave_early: {
            slave_state.fsm_state    <= slave_fsm_toggle_complete;
            slave_state.toggles.seen  <= slave_state.toggles.seen + 1;
            slave_state.toggles.early <= slave_state.toggles.early + 1;
        }
        case slave_action_slave_late: {
            slave_state.fsm_state    <= slave_fsm_toggle_complete;
            slave_state.toggles.seen <= slave_state.toggles.seen + 1;
            slave_state.toggles.late <= slave_state.toggles.late + 1;
        }
        case slave_action_unexpected_toggle: {
            slave_state.fsm_state    <= slave_fsm_toggle_complete;
            slave_state.toggles.seen <= slave_state.toggles.seen + 1;
            slave_state.toggles.unexpected <= 1;
        }
        case slave_action_not_locked: {
            slave_state.fsm_state    <= slave_fsm_idle;
            slave_state.toggles <= {*=0};
            slave_state.phase_locked <= 0;
            slave_state.locked <= 0;
        }
        case slave_action_locked: {
            slave_state.fsm_state    <= slave_fsm_idle;
            slave_state.toggles <= {*=0};
            slave_state.phase_locked <= 1;
            slave_state.locked <= slave_combs.top_value_matches;
            slave_state.request_timing <= timing_op_none;
        }
        case slave_action_locked_retard: {
            slave_state.fsm_state    <= slave_fsm_idle;
            slave_state.toggles <= {*=0};
            slave_state.phase_locked <= 1;
            slave_state.locked <= slave_combs.top_value_matches;
            slave_state.request_timing <= timing_op_retard;
        }
        case slave_action_locked_advance: {
            slave_state.fsm_state    <= slave_fsm_idle;
            slave_state.toggles <= {*=0};
            slave_state.phase_locked <= 1;
            slave_state.locked <= slave_combs.top_value_matches;
            slave_state.request_timing <= timing_op_advance;
        }
        }

        /*b Record the timer_control required */
        slave_state.timer_control.reset_counter  <= slave_sync_master_reset_counter;
        slave_state.timer_control.enable_counter <= slave_sync_master_enable_counter;
        slave_state.timer_control.lock_to_master <= slave_sync_master_lock_to_master;
        slave_state.timer_control.advance <= 0;
        slave_state.timer_control.retard  <= 0;
        if (slave_state.request_timing != timing_op_none) {
            slave_state.request_timing <= timing_op_none;
            if (slave_sync_master_lock_to_master) {
                slave_state.timer_control.advance <= (slave_state.request_timing==timing_op_advance);
                slave_state.timer_control.retard  <= (slave_state.request_timing==timing_op_retard);
            }
        }
        slave_state.synchronize_request <= slave_sync_master_synchronize_request;
        slave_state.timer_control.synchronize <= 0;
        if (!slave_sync_master_synchronize_request && slave_state.synchronize_request) { // negative edge
            slave_state.timer_control.synchronize <= 2b11;
            slave_state.timer_control.synchronize_value <= master_combs.top_value | master_combs.quarter_window;
        }
        slave_state.timer_control.block_writes            <= slave_timer_control_in.block_writes;
        slave_state.timer_control.bonus_subfraction_add   <= slave_timer_control_in.bonus_subfraction_add;
        slave_state.timer_control.bonus_subfraction_sub   <= slave_timer_control_in.bonus_subfraction_sub;
        slave_state.timer_control.fractional_adder        <= slave_timer_control_in.fractional_adder;
        slave_state.timer_control.integer_adder           <= slave_timer_control_in.integer_adder;
        slave_state.timer_control.lock_window_lsb         <= slave_timer_control_in.lock_window_lsb;

        /*b Instantiate the timer in the slave clock domain */
        clock_timer timer(clk <- slave_clk,
                          reset_n <= slave_reset_n,
                          timer_control <= slave_state.timer_control,
                          timer_value   => slave_timer_value );

        /*b Drive outputs */
        slave_timer_control_out = slave_state.timer_control;

        /*b All done */
    }

    /*b Decode window LSB - master_control.lock_window_lsb is a slow value */
    decode_window_lsb """
    Decode the @a lock_window_lsb from the @a master_timer_control, to provide
    the master and slave timer value quarter window bits, and masks
    """: {
        full_switch (master_timer_control.lock_window_lsb) {
        case timer_lock_window_lsb_6: {
            master_combs.window_bits     = master_timer_value.value[2;6];
            master_combs.top_value_mask  = (-1)<<(6+2);
            master_combs.quarter_window  = 1<<6;
            slave_combs.window_bits      = slave_timer_value.value[2;6];
        }
        case timer_lock_window_lsb_8: {
            master_combs.window_bits     = master_timer_value.value[2;8];
            master_combs.top_value_mask  = (-1)<<(8+2);
            master_combs.quarter_window  = 1<<8;
            slave_combs.window_bits      = slave_timer_value.value[2;8];
        }
        case timer_lock_window_lsb_10: {
            master_combs.window_bits     = master_timer_value.value[2;10];
            master_combs.top_value_mask  = (-1)<<(10+2);
            master_combs.quarter_window  = 1<<10;
            slave_combs.window_bits      = slave_timer_value.value[2;10];
        }
        default: { // case timer_lock_window_lsb_4: {
            master_combs.window_bits     = master_timer_value.value[2;4];
            master_combs.top_value_mask  = (-1)<<(4+2);
            master_combs.quarter_window  = 1<<4;
            slave_combs.window_bits      = slave_timer_value.value[2;4];
        }
        }
        master_combs.top_value   = master_timer_value.value & master_combs.top_value_mask;
        slave_combs.top_value    = slave_timer_value.value   & master_combs.top_value_mask;
    }
    
    /*b Logging */
    logging """
    For simulation it is useful to be able to see when the slave timer is advanced or retarded.
    This is done using simulation logging.
    """: {
        if ((slave_state.fsm_state==slave_fsm_toggle_complete) && (slave_state.toggles.seen==sync_toggle_count)) {
            log("complete",
                "master",master_timer_value.value,
                "slave",slave_timer_value.value,
                "unexpected",slave_state.toggles.unexpected,
                "early",slave_state.toggles.early,
                "late",slave_state.toggles.late,
                "diff",slave_combs.toggle_diff
                );
        }
        if (slave_state.timer_control.advance || slave_state.timer_control.retard) {
            log("adjust",
                "master",master_timer_value.value,
                "advance",slave_state.timer_control.advance,
                "slave",slave_timer_value.value,
                "m_minus_s",master_timer_value.value-slave_timer_value.value
                );
        }
    }
        
    /*b Done
     */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
